`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module priority(
input a0,a1,a2,a3,
output s0,s1
    );
    assign s0=a3|a2;
    assign s1=a3|((~a3)&(~a2)&(~a0));

endmodule
