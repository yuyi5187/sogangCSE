`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module full_subtractor(
input A,
input B,
input b,
output bn,
output D
    );
    assign D=(A^B)^b;
    assign bn=((~A)&B)|(b&(~(A^B)));
endmodule
