`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module bool_func_first_b(
input a,
input b,
input c,
output y
    );
    assign y=~((a&b)|c);
endmodule
