`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 

//////////////////////////////////////////////////////////////////////////////////


module de_morgan_first_b(
input a,
input b,
output y
    );
    assign y=(~a)&(~b);
endmodule
