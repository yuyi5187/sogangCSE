`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 

//////////////////////////////////////////////////////////////////////////////////


module bool_func_second_a(
input a,
input b,
input c,
output y

    );
    assign y=((~a)&(~b))|(~c);
endmodule
