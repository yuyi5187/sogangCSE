`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module de_morgan_second_b(
input a,
input b,
output y
    );
    assign y=(~a)|(~b);
endmodule
