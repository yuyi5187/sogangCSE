`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module encoder(
input a,
input b,
input c,
input d,
output e0,
output e1
    );
    assign e0=(a|b);
    assign e1=(a|c);
endmodule
