`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module three_input_and_gate_b(
input a,
input b,
input c,
output d,
output y
    );
    assign d=a&b;
    assign y=d&c;
endmodule
