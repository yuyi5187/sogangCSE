`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module half_subtractor(
input A,
input B,
output b,
output D
    );
    assign D=(A^B);
    assign b= (~A)&B;
endmodule
